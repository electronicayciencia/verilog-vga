//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Sat Dec 11 17:57:47 2021

module texture0_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h18C218810862188118C218C218C218C218811881188118C218C2188118C21881;
defparam prom_inst_0.INIT_RAM_01 = 256'h188108621881188118C218C218C218C218811881088318C218C218C218C218C2;
defparam prom_inst_0.INIT_RAM_02 = 256'h088318C218810883188118C218C218C208620883188108831881088318811881;
defparam prom_inst_0.INIT_RAM_03 = 256'h08621881088318810883188108831881088308621881086218C218C218C218C2;
defparam prom_inst_0.INIT_RAM_04 = 256'h1881086218C218C218C218C218C22104210421042104210418C2188118C21881;
defparam prom_inst_0.INIT_RAM_05 = 256'h18C2188118C20862188118811881086208621881188118810862188108831881;
defparam prom_inst_0.INIT_RAM_06 = 256'h18C2188118C2088318C218C2210418C218C22104210418C218C218C218C218C2;
defparam prom_inst_0.INIT_RAM_07 = 256'h188118C2188118C20862188108620862188118C2088318810862188118811881;
defparam prom_inst_0.INIT_RAM_08 = 256'h1881088318C218C218C218C221042104088318C21881088318C218C218C218C2;
defparam prom_inst_0.INIT_RAM_09 = 256'h18C218C218C218C22104210418C2210418C218C218C218C22104210418C22104;
defparam prom_inst_0.INIT_RAM_0A = 256'h21041881188118C20883210418C2210418C2188118C21881210418C2210418C2;
defparam prom_inst_0.INIT_RAM_0B = 256'h18C218C218C221042104210421042104210418C218C2210418C2210418C22104;
defparam prom_inst_0.INIT_RAM_0C = 256'h18C218C218C218C218C21881088318811881210418C218C21881088318C218C2;
defparam prom_inst_0.INIT_RAM_0D = 256'h18C2210421042104210418811881210418C22104210418C2210418C2188118C2;
defparam prom_inst_0.INIT_RAM_0E = 256'h210418C218C2088318C218C21881188118C2210418C218C218C218C218C218C2;
defparam prom_inst_0.INIT_RAM_0F = 256'h188118C221042104188118C218C218C218C2210418C22104188118C208621881;
defparam prom_inst_0.INIT_RAM_10 = 256'h08620862086218C218C218C218C2188118C21881086218C21881088318C218C2;
defparam prom_inst_0.INIT_RAM_11 = 256'h086218811881088318C218C218C218C208621881088318C218C218C218C20862;
defparam prom_inst_0.INIT_RAM_12 = 256'h086218810862188118C2210418C218C218C218C21881088318C218C2188118C2;
defparam prom_inst_0.INIT_RAM_13 = 256'h18810862188118811881188121040862188108621881188118C218C218811881;
defparam prom_inst_0.INIT_RAM_14 = 256'h1881188118811881086208621881086218812104188118811881086208621881;
defparam prom_inst_0.INIT_RAM_15 = 256'h188118C21881088318C2188108621881086218C2088318C218810862088318C2;
defparam prom_inst_0.INIT_RAM_16 = 256'h08831881088318810862086208621881210418C2210418810862086218811881;
defparam prom_inst_0.INIT_RAM_17 = 256'h188118C208621881188118C21881086218811881188118810862188118811881;
defparam prom_inst_0.INIT_RAM_18 = 256'h18C218C218C218C2188118C218C218C218C218C2210418C22104210421042104;
defparam prom_inst_0.INIT_RAM_19 = 256'h18C218C218C218C2210421042104210418C218C2188118C221042104210418C2;
defparam prom_inst_0.INIT_RAM_1A = 256'h18C218C2088318C218C2088318C2088318C218C2210421042104210421041881;
defparam prom_inst_0.INIT_RAM_1B = 256'h18C218C218C22104210418C221042104210418C218C218C2210418C218C22104;
defparam prom_inst_0.INIT_RAM_1C = 256'h210418C218C218C218C218C218C218C221042104210421042104188118C21881;
defparam prom_inst_0.INIT_RAM_1D = 256'h210418C221042104210418C218C2210418C2210418C218C2088318C218810862;
defparam prom_inst_0.INIT_RAM_1E = 256'h18812104210418C218C218C218C218C218C22104210421041881188118811881;
defparam prom_inst_0.INIT_RAM_1F = 256'h18C2210418C2210418C218C218C218C22104210418C2088318C2188108831881;
defparam prom_inst_0.INIT_RAM_20 = 256'h088318811881210418C218C2210418C218C2188108621881086218C218C218C2;
defparam prom_inst_0.INIT_RAM_21 = 256'h188118811881086218C2088318C218810862086218C21881188118C2188118C2;
defparam prom_inst_0.INIT_RAM_22 = 256'h188118C20862188118C218C218C21881088318811881086218C218C218C218C2;
defparam prom_inst_0.INIT_RAM_23 = 256'h1881086218811881188118C2188118C2188118810862188108831881088318C2;
defparam prom_inst_0.INIT_RAM_24 = 256'h088318C218C218C20862188108620862086218811881188118C2088318C21881;
defparam prom_inst_0.INIT_RAM_25 = 256'h210421042104210418C218C2088318C2210421042104210418C218C218811881;
defparam prom_inst_0.INIT_RAM_26 = 256'h18C218C2088318810862188108620862210418C218C2188118C2188118811881;
defparam prom_inst_0.INIT_RAM_27 = 256'h210418C218C2210418C218C218C218C2210418C218812104210418C218810883;
defparam prom_inst_0.INIT_RAM_28 = 256'h18C218C218C218C2210421042104210418C218C218C2210418C22104210418C2;
defparam prom_inst_0.INIT_RAM_29 = 256'h18C218C21881086218C2088318C218C218C218C218C218C2210418C221042104;
defparam prom_inst_0.INIT_RAM_2A = 256'h18C218C218C2210418C218C22104210418C218C218C218C2210418C218C218C2;
defparam prom_inst_0.INIT_RAM_2B = 256'h18C218C208621881188118C218C218C218C218C21881088318C218C2210418C2;
defparam prom_inst_0.INIT_RAM_2C = 256'h18C218C218C218C2088318C21881088318C218C218C218C21881088318811881;
defparam prom_inst_0.INIT_RAM_2D = 256'h18C218C218810862086208620862086218C218C2188118C20883188118810883;
defparam prom_inst_0.INIT_RAM_2E = 256'h188118C218C218C21881188118811881188118C218C208621881188108831881;
defparam prom_inst_0.INIT_RAM_2F = 256'h18C2188118C21881086218810862086218C218C218C218811881188108831881;
defparam prom_inst_0.INIT_RAM_30 = 256'h08620862188118811881210418C2086218811881086208620862188118C21881;
defparam prom_inst_0.INIT_RAM_31 = 256'h18810862188118C221042104210418C218C218C20883210418C218C218C20862;
defparam prom_inst_0.INIT_RAM_32 = 256'h00211881188118812104210418C221041881086208620862188118C2188118C2;
defparam prom_inst_0.INIT_RAM_33 = 256'h1881188118C218C218C2210421042104210418C218C218C218C2210418C218C2;
defparam prom_inst_0.INIT_RAM_34 = 256'h1881088318C218C218C218C2210418C22104210418C22104210418C218C218C2;
defparam prom_inst_0.INIT_RAM_35 = 256'h2104210418C2210418C218C218C2210418C2210418C218C2088318C200210862;
defparam prom_inst_0.INIT_RAM_36 = 256'h18C21881088318C218C218C218C2210418C221042104210418C218C218C218C2;
defparam prom_inst_0.INIT_RAM_37 = 256'h2104210421041881088318C2088318C21881210418C218C218C2086208621881;
defparam prom_inst_0.INIT_RAM_38 = 256'h210418C218C218C218C22104210418C218C218C2188118C218C2210421042104;
defparam prom_inst_0.INIT_RAM_39 = 256'h18811881086218C2188118C218C218C2088318810883188118C218C221041881;
defparam prom_inst_0.INIT_RAM_3A = 256'h18C2210418C218C218C218C218C218C2088318C218C20883210418C221042104;
defparam prom_inst_0.INIT_RAM_3B = 256'h188108831881188118C218C218C20883188118C2188118C21881210421042104;
defparam prom_inst_0.INIT_RAM_3C = 256'h2104210418C22104088318810883188118C218C218C218811881188118811881;
defparam prom_inst_0.INIT_RAM_3D = 256'h21042104210418810883188118C21881188118C218C218C218C2188118C218C2;
defparam prom_inst_0.INIT_RAM_3E = 256'h18812104210418811881188118811881188118C218C218C21881086218811881;
defparam prom_inst_0.INIT_RAM_3F = 256'h18C218C218C218C21881188118811881210418C218C2188108831881188118C2;

endmodule //texture0_rom
