//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.03
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Wed Nov 01 18:10:35 2023

module charbuf_color_64x32 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [10:0] ada;
input [15:0] din;
input [10:0] adb;

wire [23:0] sdpb_inst_0_dout_w;
wire [23:0] sdpb_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[23:0],dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 8;
defparam sdpb_inst_0.BIT_WIDTH_1 = 8;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDC9;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h00000000BBCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCD;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h342044434C202020206F6D656420414756206B31206F6E614E20676E615420BA;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h00000000BA203731783036202074786574203631783820202020323732783038;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hC4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C7;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h00000000B6C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h20202020202020202020202020202020202020202020202020202020202020BA;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h00000000BA202020202020202020202020202020202020202020202020202020;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h36353433323130202020202046454443424139383736353433323130202020BA;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h00000000BA202073726F6C6F4320746962382020202020464544434241393837;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h8685848382818038202020200F0E0D0C0B0A09080706050403020100302020BA;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h00000000BA20206161DBDB3820206161DBDB30202020208F8E8D8C8B8A898887;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h9695949392919039202020201F1E1D1C1B1A19181716151413121110312020BA;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h00000000BA20206161DBDB3920206161DBDB31202020209F9E9D9C9B9A999897;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hA6A5A4A3A2A1A041202020202F2E2D2C2B2A29282726252423222120322020BA;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h00000000BA20206161DBDB3031206161DBDB3220202020AFAEADACABAAA9A8A7;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hB6B5B4B3B2B1B042202020203F3E3D3C3B3A39383736353433323130332020BA;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h00000000BA20206161DBDB3131206161DBDB3320202020BFBEBDBCBBBAB9B8B7;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hC6C5C4C3C2C1C043202020204F4E4D4C4B4A49484746454443424140342020BA;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h00000000BA20206161DBDB3231206161DBDB3420202020CFCECDCCCBCAC9C8C7;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hD6D5D4D3D2D1D044202020205F5E5D5C5B5A59585756555453525150352020BA;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h00000000BA20206161DBDB3331206161DBDB3520202020DFDEDDDCDBDAD9D8D7;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hE6E5E4E3E2E1E045202020206F6E6D6C6B6A69686766656463626160362020BA;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h00000000BA20206161DBDB3431206161DBDB3620202020EFEEEDECEBEAE9E8E7;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hF6F5F4F3F2F1F046202020207F7E7D7C7B7A79787776757473727170372020BA;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h00000000BA20206161DBDB3531206161DBDB3720202020FFFEFDFCFBFAF9F8F7;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h20202020202020202020202020202020202020202020202020202020202020BA;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h00000000BA202020202020202020202020202020202020202020202020202020;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hC4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C7;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h00000000B6C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h202020206169636E6569432079206163696EA2727463656C4520676F6C4220BA;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h00000000BA20333230322F31312F313020202020202020202020202020202020;
defparam sdpb_inst_0.INIT_RAM_20 = 256'hCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDC8;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h00000000BCCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCD;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[23:0],dout[15:8]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:8]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 8;
defparam sdpb_inst_1.BIT_WIDTH_1 = 8;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h0000000001010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h0202020202020202020202020202020202020202020202020202020202020001;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h0000000001000202020202020202020202020202020202020202020202020202;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h0000000001010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000001;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h0000000001000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h0F0F0F0F0F0F0F00000000000F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F00000001;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h000000000100000F0F0F0F0F0F0F0F0F0F0F00000000000F0F0F0F0F0F0F0F0F;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h00000000010000088008080F0F00000000000F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h00000000010000099009090F0F00011001010F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h000000000100000AA00A0A0F0F00022002020F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h000000000100000BB00B0B0F0F00033003030F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h000000000100000CC00C0C0F0F00044004040F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h000000000100000DD00D0D0F0F00055005050F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h000000000100000EE00E0E0F0F00066006060F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h070707070707070F00000000070707070707070707070707070707070F000001;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h000000000100000FF00F0F0F0F00077007070F00000000070707070707070707;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000001;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h0000000001000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0000000001010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h0303030303030303030303030303030303030303030303030303030303030001;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h0000000001000303030303030303030303030303030303030303030303030303;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h0000000001010101010101010101010101010101010101010101010101010101;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //charbuf_color_64x32
