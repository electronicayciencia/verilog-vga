//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Wed Dec 15 18:38:42 2021

module charbuf_mono_64x64 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [11:0] ada;
input [7:0] din;
input [11:0] adb;

wire [27:0] sdpb_inst_0_dout_w;
wire [27:0] sdpb_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[27:0],dout[3:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 4;
defparam sdpb_inst_0.BIT_WIDTH_1 = 4;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h00003210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA98;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h0000FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA987654;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h0000BA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h000076543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDC;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[27:0],dout[7:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 4;
defparam sdpb_inst_1.BIT_WIDTH_1 = 4;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h3333333333333333222222222222222211111111111111110000000000000000;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h3333777777776666666666666666555555555555555544444444444444443333;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h3333BBBBAAAAAAAAAAAAAAAA9999999999999999888888888888888877777777;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h3333EEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCBBBBBBBBBBBB;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h333322222222222211111111111111110000000000000000FFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h3333666666665555555555555555444444444444444433333333333333332222;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h3333AAAA99999999999999998888888888888888777777777777777766666666;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h3333DDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAA;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h33331111111111110000000000000000FFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEE;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h3333555555554444444444444444333333333333333322222222222222221111;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h3333999988888888888888887777777777777777666666666666666655555555;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h3333CCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h3333000000000000FFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDD;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h3333444444443333333333333333222222222222222211111111111111110000;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h3333888877777777777777776666666666666666555555555555555544444444;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h3333BBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA9999999999999999888888888888;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h3333FFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCC;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h333333333333222222222222222211111111111111110000000000000000FFFF;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h3333777766666666666666665555555555555555444444444444444433333333;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h3333AAAAAAAAAAAAAAAA99999999999999998888888888888888777777777777;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h3333EEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBB;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h33332222222211111111111111110000000000000000FFFFFFFFFFFFFFFFEEEE;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h3333666655555555555555554444444444444444333333333333333322222222;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h3333999999999999999988888888888888887777777777777777666666666666;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h3333DDDDDDDDDDDDCCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h3333111111110000000000000000FFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDD;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h3333555544444444444444443333333333333333222222222222222211111111;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h3333888888888888888877777777777777776666666666666666555555555555;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h3333CCCCCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA9999999999999999;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h333300000000FFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCC;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h3333444433333333333333332222222222222222111111111111111100000000;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h3333777777777777777766666666666666665555555555555555444444444444;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h3333BBBBBBBBBBBBAAAAAAAAAAAAAAAA99999999999999998888888888888888;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h3333FFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCBBBB;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h3333333333333333333333333333333333333333333333333333333333333333;

endmodule //charbuf_mono_64x64
