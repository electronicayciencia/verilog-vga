//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.03
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Wed Nov 15 21:33:16 2023

module vram_m64x32 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [10:0] ada;
input [7:0] dina;
input [10:0] adb;
input [7:0] dinb;

wire [7:0] dpb_inst_0_douta_w;
wire [7:0] dpb_inst_0_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[7:0],douta[7:0]}),
    .DOB({dpb_inst_0_doutb_w[7:0],doutb[7:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b01;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 8;
defparam dpb_inst_0.BIT_WIDTH_1 = 8;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h797563206564202C6168636E614D20616C20656420726167756C206E75206E45;
defparam dpb_inst_0.INIT_RAM_01 = 256'h20202020202D726164726F6361206F7265697571206F6E206572626D6F6E206F;
defparam dpb_inst_0.INIT_RAM_02 = 256'h61A176697620657571206F706D656974206F6863756D206168206F6E202C656D;
defparam dpb_inst_0.INIT_RAM_03 = 256'h2020202020617A6E616C20656420736F6C206564206F676C61646968206E7520;
defparam dpb_inst_0.INIT_RAM_04 = 256'h6F72202C61756769746E6120616772616461202C6F72656C6C69747361206E65;
defparam dpb_inst_0.INIT_RAM_05 = 256'h20202020202E726F646572726F63206F676C61672079206F63616C66206EA163;
defparam dpb_inst_0.INIT_RAM_06 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_07 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_08 = 256'h61632065757120616361762073A06D206F676C6120656420616C6C6F20616E55;
defparam dpb_inst_0.INIT_RAM_09 = 256'h20202020202D6F6E2073A06D2073616C206EA26369706C6173202C6F72656E72;
defparam dpb_inst_0.INIT_RAM_0A = 256'hA07320736F6C20736F746E617262657571207920736F6C657564202C73656863;
defparam dpb_inst_0.INIT_RAM_0B = 256'h202020202C73656E7265697620736F6C2073616A65746E616C202C736F646162;
defparam dpb_inst_0.INIT_RAM_0C = 256'h20736F6C2061727564696461A461206564206F6E696D6F6C6170206EA3676C61;
defparam dpb_inst_0.INIT_RAM_0D = 256'h20202020736572742073616C206E61A16D75736E6F63202C736F676E696D6F64;
defparam dpb_inst_0.INIT_RAM_0E = 256'h206F74736572206C45202E61646E656963616820757320656420736574726170;
defparam dpb_inst_0.INIT_RAM_0F = 256'h20202020202D6576206564206F796173206E61A1756C636E6F6320616C6C6564;
defparam dpb_inst_0.INIT_RAM_10 = 256'h616C2061726170206F64756C6C65762065642073617A6C6163202C657472616C;
defparam dpb_inst_0.INIT_RAM_11 = 256'h20202020736F6C6675746E617020737573206E6F63202C736174736569662073;
defparam dpb_inst_0.INIT_RAM_12 = 256'h6572746E65206564207361A16420736F6C2079202C6F6D73656D206F6C206564;
defparam dpb_inst_0.INIT_RAM_13 = 256'h20202020202020207573206E6F6320616261726E6F6820657320616E616D6573;
defparam dpb_inst_0.INIT_RAM_14 = 256'h2020202020202020202E6F6E69662073A06D206F6C20656420A1726F6C6C6576;
defparam dpb_inst_0.INIT_RAM_15 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_16 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_17 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_18 = 256'h7361702065757120616D6120616E752061736163207573206E652061A16E6554;
defparam dpb_inst_0.INIT_RAM_19 = 256'h20202020202020616E7520792061746E657261756320736F6C20656420616261;
defparam dpb_inst_0.INIT_RAM_1A = 256'h69657620736F6C20612061626167656C6C206F6E2065757120616E6972626F73;
defparam dpb_inst_0.INIT_RAM_1B = 256'h2020202020202079206F706D6163206564206F7A6F6D206E752079202C65746E;
defparam dpb_inst_0.INIT_RAM_1C = 256'h6EA1636F72206C65206162616C6C69736E6520A173612065757120617A616C70;
defparam dpb_inst_0.INIT_RAM_1D = 256'h202020202020202E6172656461646F7020616C206162616D6F74206F6D6F6320;
defparam dpb_inst_0.INIT_RAM_1E = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_1F = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_20 = 256'h6C61646968206F72747365756E206564206461646520616C2061626173697246;
defparam dpb_inst_0.INIT_RAM_21 = 256'h2020202020202E736FA4612061746E6575636E696320736F6C206E6F63206F67;
defparam dpb_inst_0.INIT_RAM_22 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_23 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_24 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_25 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_26 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_27 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_28 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_29 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_2A = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_2B = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_2C = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_2D = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_2E = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_2F = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_30 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_31 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_32 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_33 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_34 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_35 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_36 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_37 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_38 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_39 = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_3A = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_3B = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_3C = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_3D = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_3E = 256'h2020202020202020202020202020202020202020202020202020202020202020;
defparam dpb_inst_0.INIT_RAM_3F = 256'h2020202020202020202020202020202020202020202020202020202020202020;

endmodule //vram_m64x32
