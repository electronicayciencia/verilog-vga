//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.03
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Mon Oct 09 16:09:10 2023

module charbuf_mono_64x64 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [11:0] ada;
input [7:0] din;
input [11:0] adb;

wire [27:0] sdpb_inst_0_dout_w;
wire [27:0] sdpb_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[27:0],dout[3:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 4;
defparam sdpb_inst_0.BIT_WIDTH_1 = 4;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h00000000000000A5EFD94E5740F405E9E03532560CF74025401830C34E5D1D21;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h000007E99130C87980EF0050541E52704E180584045391201C944104E91304E1;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000541E52704E180984039840335C20C42FC0F2;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h00000003749209E940F40359D5E505E98407FC2043591D05F840490849704184;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h000000000000000000000000000000000000000000000000002E9325D09840E9;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h000000005840EF05043156049405C0F50058404E10CE9270494042FC058404E1;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h0000003E1457E12F04E10C3596F83E104E10C021304E10C384FC304E10C32D1C;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h0000000000EEE58305721C04E10341204952604E103C152530C4316B152204E1;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000A7E99130C5B103042FC058404E1;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000E9009CF80584045F05B1405F8404C1830432962;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000552840F404E5F305F8404C1830E584;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000335C0FE052FD0FE;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h00000000000000000000004E5F304C18305F840252D5E058405204C183055284;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h0000000000000000000552840520CC18307E94E5F3058406F0252D5E058404E1;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000004E5F304FE05F8404C183025F6;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h000000000000000000000000000000000000000F7405F8404E5F3025849502FE;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h00000000000000000000000552840F404553F200E58405F840418407E9405385;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000045F04879203905696;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h000000045831520520C252D5E042984058407E9520C552840252D5E0584053EF;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h00000034217F4083F94E106F0541E52704E1809CF8098405F84043522FC0E584;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h000000002490665E30CC1830C4879309D0E90948751E07E9520CF870C5F60984;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h000000000000000000000000000000000000000000000000000000000000E5D1;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[27:0],dout[7:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 4;
defparam sdpb_inst_1.BIT_WIDTH_1 = 4;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h2222222222222236662776677267266662767767226772767766622776666674;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h2222266676722666626627726666674266662667266766726667742766652664;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h2222222222222222222222222222666667426666276527667277666226764242;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h2222222727662766526727666666266665276662776766276652762676727665;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h2222222222222222222222222222222222222222222222222222767662765264;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h2222222266726677277666266626676672667266622667626662676426672664;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h2222227667766676266622766766666266622776626662276766726662276666;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h2222222222222766266766266627766276776266627666766227766666762666;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h2222222222222222222222222222222222222366676722666772676426672664;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h2222222222222222222222222665276642667277626667276672766672777642;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h2222222222222222222222222222222222667672672767662766727666726665;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h2222222222222222222222222222222222222222222222222776626626766264;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h2222222222222222222222767662766672766727666762667266276667266765;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h2222222222222222222667672662666672666767662667266276667626672664;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h2222222222222222222222222222222222222227676627662766727666727764;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h2222222222222222222222222222222222222226772766727676627667662764;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h2222222222222222222222266765267266666772666727667276672666776674;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h2222222222222222222222222222222222222222222222277627666727626764;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h2222222666666726622766676267667266726666622667672766676266726664;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h2222227676767266667642662666667426664276642765276672776666626665;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h2222222227626676726666722766672742662776676626666622667226662765;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h2222222222222222222222222222222222222222222222222222222222226664;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h2222222222222222222222222222222222222222222222222222222222222222;

endmodule //charbuf_mono_64x64
