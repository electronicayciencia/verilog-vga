//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Sat Dec 11 17:45:11 2021

module texture1_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h188118811881188118C218C218C218C218811881188118811881188118C218C2;
defparam prom_inst_0.INIT_RAM_01 = 256'h18C218C218C218C218C218C218C2188118811881188118811881188118811881;
defparam prom_inst_0.INIT_RAM_02 = 256'h28C23964396439643964396441844184418441844184418439643964396418C2;
defparam prom_inst_0.INIT_RAM_03 = 256'h28C228C2396428C24184418441844184418441843964396428C228C228C21881;
defparam prom_inst_0.INIT_RAM_04 = 256'h20A528C228C228C228C228C228C228C220A528C228C220A528C228C228C218C2;
defparam prom_inst_0.INIT_RAM_05 = 256'h18C228C228C228C228C228C220A528C228C220A528C228C228C228C228C218C2;
defparam prom_inst_0.INIT_RAM_06 = 256'h280028C220A528C228C220A5404020A5412228C228C2412220A528C228C228C2;
defparam prom_inst_0.INIT_RAM_07 = 256'h18C228C220A528C220A528C2404020A5412228C228C220A528C228C2396418C2;
defparam prom_inst_0.INIT_RAM_08 = 256'h20A528C220A5404020A5412220A5412220A558A220A528C228C228C228C218C2;
defparam prom_inst_0.INIT_RAM_09 = 256'h18C228C228C228C228C228C220A5412220A528C228C228C228C228C228C21881;
defparam prom_inst_0.INIT_RAM_0A = 256'h18C228C228C228C228C228C228C228C228C220A528C228C220A5412228C228C2;
defparam prom_inst_0.INIT_RAM_0B = 256'h18C228C220A5412220A5412228C228C228C220A528C228C220A528C228C218C2;
defparam prom_inst_0.INIT_RAM_0C = 256'h1881188118C220A528C220A528C220A528C228C228C228C2412220A528C218C2;
defparam prom_inst_0.INIT_RAM_0D = 256'h18C228C228C228C228C220A528C220A528C228C220A528C228C228C239641881;
defparam prom_inst_0.INIT_RAM_0E = 256'h18811881188118C228C228C228C228C218C218C218C218C228C228C228C228C2;
defparam prom_inst_0.INIT_RAM_0F = 256'h18C218C218C218C228C228C228C228C228C218C228C228C228C228C228C218C2;
defparam prom_inst_0.INIT_RAM_10 = 256'h28001881188118811881188118811881188118C2280018C2188118C218C218C2;
defparam prom_inst_0.INIT_RAM_11 = 256'h18C2280018811881188118811881188108832800088328000883188118810883;
defparam prom_inst_0.INIT_RAM_12 = 256'h39644184418441844184418441844184418441843964188128C228C228C23964;
defparam prom_inst_0.INIT_RAM_13 = 256'h28C228C228C228C228C228C23964396439643964396418813964396439643964;
defparam prom_inst_0.INIT_RAM_14 = 256'h20A528C220A528C220A528C220A528C220A528C228C228C220A528C228C228C2;
defparam prom_inst_0.INIT_RAM_15 = 256'h28C228C220A5396428C220A528C228C228C228C2396420A528C228C220A54040;
defparam prom_inst_0.INIT_RAM_16 = 256'h28C228C228C258A220A54040396428C228C228C228C218C218C228C228C220A5;
defparam prom_inst_0.INIT_RAM_17 = 256'h210428C228C228C228C228C228C220A528C228C23964280028C228C228C228C2;
defparam prom_inst_0.INIT_RAM_18 = 256'h28C220A528C220A5412220A528C228C220A528C228C21881280020A528C228C2;
defparam prom_inst_0.INIT_RAM_19 = 256'h28C228C220A528C228C220A528C228C228C228C2418428C220A528C228C220A5;
defparam prom_inst_0.INIT_RAM_1A = 256'h28C228C228C228C228C228C228C228C228C228C228C218C218C228C228C228C2;
defparam prom_inst_0.INIT_RAM_1B = 256'h18C228C228C228C228C228C228C220A528C228C228C228C228C228C228C228C2;
defparam prom_inst_0.INIT_RAM_1C = 256'h28C228C220A558A220A5412220A528C220A528C228C2188118C218C218C228C2;
defparam prom_inst_0.INIT_RAM_1D = 256'h28C220A528C228C228C218C218C228C228C228C228C218C218C220A528C220A5;
defparam prom_inst_0.INIT_RAM_1E = 256'h18C228C218C228C228C218C228C228C228C228C228C218C218C2280018C218C2;
defparam prom_inst_0.INIT_RAM_1F = 256'h18C218C228C220A528C218C218C228C218C228C228C218C21881188118C228C2;
defparam prom_inst_0.INIT_RAM_20 = 256'h18C2188118C2188118C2188118811881188118811881188118C218C218C218C2;
defparam prom_inst_0.INIT_RAM_21 = 256'h18C218C218C218C2280020A5280018C218C218C228C218C2280018C218811881;
defparam prom_inst_0.INIT_RAM_22 = 256'h3964396439643964396439643964188128C228C2396428C228C2396428C228C2;
defparam prom_inst_0.INIT_RAM_23 = 256'h28C228C2412228C2396428C228C218C228C228C228C2396428C228C239641881;
defparam prom_inst_0.INIT_RAM_24 = 256'h28C228C228C228C228C228C228C228C220A528C228C220A528C228C228C218C2;
defparam prom_inst_0.INIT_RAM_25 = 256'h28C228C220A528C220A528C228C218C228C220A528C228C228C228C2396420A5;
defparam prom_inst_0.INIT_RAM_26 = 256'h280020A528C220A528C228C228C228C228C228C228C228C228C220A5412218C2;
defparam prom_inst_0.INIT_RAM_27 = 256'h210428C228C228C228C228C228C2188128C228C228C220A528C228C2396418C2;
defparam prom_inst_0.INIT_RAM_28 = 256'h20A528C228C228C228C228C228C218C220A528C228C220A528C228C228C218C2;
defparam prom_inst_0.INIT_RAM_29 = 256'h28C228C228C220A528C228C228C2188128C220A528C228C228C228C2396428C2;
defparam prom_inst_0.INIT_RAM_2A = 256'h280028C220A528C228C220A528C228C228C228C228C228C228C228C2396418C2;
defparam prom_inst_0.INIT_RAM_2B = 256'h210428C228C228C228C220A528C2188118C228C228C228C220A528C228C218C2;
defparam prom_inst_0.INIT_RAM_2C = 256'h20A528C228C228C228C228C228C218C220A528C228C218C228C218C228C218C2;
defparam prom_inst_0.INIT_RAM_2D = 256'h28C228C220A528C228C228C228C2188118C228C228C228C228C228C228C218C2;
defparam prom_inst_0.INIT_RAM_2E = 256'h18C218C228C228C218C228C228C228C228C228C218C218C218C218C228C218C2;
defparam prom_inst_0.INIT_RAM_2F = 256'h18C228C228C228C220A528C228C218C218C218C218C228C218C218C228C218C2;
defparam prom_inst_0.INIT_RAM_30 = 256'h1881188118C218C2188118811881188118811881188118812800188118C218C2;
defparam prom_inst_0.INIT_RAM_31 = 256'h18C218C218C218C2188118C218C218C21881188118C218C2188118C218811881;
defparam prom_inst_0.INIT_RAM_32 = 256'h28C2396428C2396428C239643964396441844184418439643964396439641881;
defparam prom_inst_0.INIT_RAM_33 = 256'h28C2418441844184418441844184418441844184418439643964396428C21881;
defparam prom_inst_0.INIT_RAM_34 = 256'h28C228C228C228C228C228C228C228C220A528C228C220A528C228C228C228C2;
defparam prom_inst_0.INIT_RAM_35 = 256'h18C228C220A528C220A528C220A528C220A528C220A528C228C228C228C218C2;
defparam prom_inst_0.INIT_RAM_36 = 256'h28C220A528C220A528C220A528C228C228C228C228C258A220A528C258A220A5;
defparam prom_inst_0.INIT_RAM_37 = 256'h28C228C228C228C228C228C228C228C228C228C228C228C220A528C228C218C2;
defparam prom_inst_0.INIT_RAM_38 = 256'h28C228C228C228C228C228C228C220A5404020A528C220A5412220A528C218C2;
defparam prom_inst_0.INIT_RAM_39 = 256'h18C220A528C228C220A528C228C220A528C228C220A528C228C228C228C218C2;
defparam prom_inst_0.INIT_RAM_3A = 256'h28C220A528C228C220A558A220A528C228C228C228C228C228C228C2396418C2;
defparam prom_inst_0.INIT_RAM_3B = 256'h18C228C228C228C228C228C228C228C228C228C228C228C228C2396428C218C2;
defparam prom_inst_0.INIT_RAM_3C = 256'h18C2280028C228C228C220A528C228C228C220A528C228C220A528C228C218C2;
defparam prom_inst_0.INIT_RAM_3D = 256'h18C228C228C220A528C228C228C220A528C220A528C228C220A528C228C21881;
defparam prom_inst_0.INIT_RAM_3E = 256'h1881188118C2188118C228C228C228C218C228C218C228C228C228C228C218C2;
defparam prom_inst_0.INIT_RAM_3F = 256'h18C218C218C218C21881188118C218C218C218C228C228C218C218C228C218C2;

endmodule //texture1_rom
