//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Fri Dec 03 14:38:56 2021

module rom_4c (dout, clk, oce, ce, reset, ad);

output [1:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [1:1] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [1:1] prom_inst_3_dout;
wire dff_q_0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_1.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000800000000000000000000000000000070000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_0C = 256'h00008000000000000000000000000000000703FC000000000000000000000001;
defparam prom_inst_0.INIT_RAM_0D = 256'h00008000000000000000000000000000000707FC000000000000000000000001;
defparam prom_inst_0.INIT_RAM_0E = 256'h000080000000000000000000000000000007070C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_0F = 256'h00008000000000000000000000003F807E07060C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_10 = 256'h00008000000000000000000000003FC0FF07060C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_11 = 256'h000080000000000000000000000039E0E787070C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_12 = 256'h000080000000000000000000000030E1C38703FC000000000000000000000001;
defparam prom_inst_0.INIT_RAM_13 = 256'h00008000000000000000000000003061C1870FFC000000000000000000000001;
defparam prom_inst_0.INIT_RAM_14 = 256'h00008000000000000000000000003061C1870E0C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_15 = 256'h00008000000000000000000000003061C1871C0C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_16 = 256'h00008000000000000000000000003061C3871C0C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_17 = 256'h000080000000000000000000000039E0E7870F0C000000000000000000000001;
defparam prom_inst_0.INIT_RAM_18 = 256'h00008000000000000000000000003FC0FF070FFC000000000000000000000001;
defparam prom_inst_0.INIT_RAM_19 = 256'h00008000000000000000000000003F807E0703FC000000000000000000000001;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000800000000000000000000000300000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000800000000000000000000000380000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_1C = 256'h00008000000000000000000000001FC000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_1D = 256'h00008000000000000000000000000FC000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_22 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_26 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_28 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_29 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_2A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_2C = 256'h0000800000000000000000000000000000000000000038000000000000380001;
defparam prom_inst_0.INIT_RAM_2D = 256'h00008000380000000000E000000000000000001C00001C000038000000387FC1;
defparam prom_inst_0.INIT_RAM_2E = 256'h00008000380000000000E000000000000000001C00000C000038000000387FC1;
defparam prom_inst_0.INIT_RAM_2F = 256'h00008000000000000000000000000000000000000000000000380000003800C1;
defparam prom_inst_0.INIT_RAM_30 = 256'h000083F8387E01FE0FC0E1F8001C1C001FC1F81C0FF03F07F1FC7E03F03800C1;
defparam prom_inst_0.INIT_RAM_31 = 256'h000087F838FF03FE1FE0E3FC000C18003FC3FC1C1FF07F8FF1FCFF07F83800C1;
defparam prom_inst_0.INIT_RAM_32 = 256'h0000870038E783BE1CF0E39E000E380038039E1C1DF073C0F038E7873C387FC1;
defparam prom_inst_0.INIT_RAM_33 = 256'h000086003803870E3830E00E000E300030000E1C3870E1C07038038E0C387FC1;
defparam prom_inst_0.INIT_RAM_34 = 256'h000087F03801870E3FF0E006000670003F80061C3870E0C07038018FFC3800C1;
defparam prom_inst_0.INIT_RAM_35 = 256'h000087FC3801870E3FF0E006000770003FE0061C3870E0C07038018FFC3800C1;
defparam prom_inst_0.INIT_RAM_36 = 256'h0000863C3801870E0030E0060003600031E0061C3870E0C0703801800C3800C1;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000860C3803870E0070E00E0003E00030600E1C3870E1C0703803801C3800C1;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000879C38E7870E38F0E39E0003C0003CE39E1C387073C07030E78E3C3800C1;
defparam prom_inst_0.INIT_RAM_39 = 256'h000087FC38FF070E3FE0E3FC0001C0003FE3FC1C38707F8071F0FF0FF8387FC1;
defparam prom_inst_0.INIT_RAM_3A = 256'h000086F8387E070E1FC0E1F80001C00037C1F81C38703F0071E07E07F0387FC1;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000800000000000000000000000C00000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000800000000000000000000000E00000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000800000000000000000000000E00000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000800000000000000000000000600000000000000000000000000000000001;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000800000000000000000000000000000000000000000000000000000000001;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_04 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_0A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_0C = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_0E = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_0F = 256'h00008000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000001;
defparam prom_inst_1.INIT_RAM_10 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_11 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_12 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_13 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_14 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_15 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_16 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_17 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_18 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_19 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_1A = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_1B = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_1C = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_1D = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_1E = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_1F = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_20 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_21 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_22 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_23 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_24 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_25 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_26 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_27 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_28 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_29 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_2A = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_2B = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_2C = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_2D = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_2E = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_2F = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_30 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFC000000010000000000001;
defparam prom_inst_1.INIT_RAM_31 = 256'h00008000000000001FFFFFFFFC00000001FFFFFFFFFFFFFFFFF0000000000001;
defparam prom_inst_1.INIT_RAM_32 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_33 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_34 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_35 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_36 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_37 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_01 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_02 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_03 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_04 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_05 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_06 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_07 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_08 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_09 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_0A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_0B = 256'h0000800000000000000000000000000000060000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_0C = 256'h00008000000000000000000000000000000603FC000000000000000000000001;
defparam prom_inst_2.INIT_RAM_0D = 256'h00008000000000000000000000000000000607FC000000000000000000000001;
defparam prom_inst_2.INIT_RAM_0E = 256'h000080000000000000000000000000000006070C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_0F = 256'h00008000000000000000000000003F003E06060C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_10 = 256'h00008000000000000000000000003FC07F06060C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_11 = 256'h000080000000000000000000000030C0E306030C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_12 = 256'h00008000000000000000000000003060C18603FC000000000000000000000001;
defparam prom_inst_2.INIT_RAM_13 = 256'h00008000000000000000000000003061818607FC000000000000000000000001;
defparam prom_inst_2.INIT_RAM_14 = 256'h0000800000000000000000000000306181860E0C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_15 = 256'h0000800000000000000000000000306181860C0C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_16 = 256'h00008000000000000000000000003060C1860C0C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_17 = 256'h000080000000000000000000000038E0E3060E0C000000000000000000000001;
defparam prom_inst_2.INIT_RAM_18 = 256'h00008000000000000000000000003FC07F0607FC000000000000000000000001;
defparam prom_inst_2.INIT_RAM_19 = 256'h000080000000000000000000000037803E0603FC000000000000000000000001;
defparam prom_inst_2.INIT_RAM_1A = 256'h0000800000000000000000000000300000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000800000000000000000000000380000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_1C = 256'h00008000000000000000000000001FC000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_1D = 256'h00008000000000000000000000000FC000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_1E = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_1F = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_20 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_21 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_22 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_23 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_24 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_25 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_26 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_27 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_28 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_29 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_2A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_2B = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_2C = 256'h0000800000000000000000000000000000000000000018000000000000300001;
defparam prom_inst_2.INIT_RAM_2D = 256'h00008000300000000000C000000000000000001800000C000030000000307FC1;
defparam prom_inst_2.INIT_RAM_2E = 256'h00008000300000000000C000000000000000001800000C000030000000307FC1;
defparam prom_inst_2.INIT_RAM_2F = 256'h00008000000000000000000000000000000000000000000000300000003000C1;
defparam prom_inst_2.INIT_RAM_30 = 256'h000081F8307C01EC0780C1F0001818000FC1F0180F601F0761FC7C01E03000C1;
defparam prom_inst_2.INIT_RAM_31 = 256'h000083F8307F03FC0FE0C1FC000C18001FC1FC181FE03F87E1FC7F03F83000C1;
defparam prom_inst_2.INIT_RAM_32 = 256'h000087003043031C1860C10C000C380038010C1818E07180E030430618307FC1;
defparam prom_inst_2.INIT_RAM_33 = 256'h000086003001830C1830C0060006300030000618186060C0603001860C307FC1;
defparam prom_inst_2.INIT_RAM_34 = 256'h000087F03001820C1FF0C006000630003F8006181060C0C060300187FC3000C1;
defparam prom_inst_2.INIT_RAM_35 = 256'h000087F83001820C1FF0C006000760003FC006181060C0C060300187FC3000C1;
defparam prom_inst_2.INIT_RAM_36 = 256'h0000861C3001820C0030C0060003600030E006181060C0C0603001800C3000C1;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000860C3001820C0030C0060003E00030600618106060C0603001800C3000C1;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000870C3043020C1060C10C0001C00038610C181060718060304304183000C1;
defparam prom_inst_2.INIT_RAM_39 = 256'h000087FC307F020C1FE0C1FC0001C0003FE1FC1810603F8061F07F07F8307FC1;
defparam prom_inst_2.INIT_RAM_3A = 256'h000086F8307E020C0F80C1F80001C00037C1F81810601F0061E07E03E0307FC1;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000800000000000000000000000C00000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000800000000000000000000000C00000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000800000000000000000000000600000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000800000000000000000000000600000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000800000000000000000000000000000000000000000000000000000000001;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_01 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_02 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_03 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_04 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_05 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_06 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_07 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_08 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_09 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_0A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_0B = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_0C = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_0D = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_0E = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_0F = 256'h00008000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000001;
defparam prom_inst_3.INIT_RAM_10 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_11 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_12 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_13 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_14 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_15 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_16 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_17 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_18 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_19 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_1A = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_1B = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_1C = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_1D = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_1E = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_1F = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_20 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_21 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_22 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_23 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_24 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_25 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_26 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_27 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_28 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_29 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_2A = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_2B = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_2C = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_2D = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_2E = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_2F = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_30 = 256'h00008000000000001FFFFFFFFFFFFFFFFF000000004000000010000000000001;
defparam prom_inst_3.INIT_RAM_31 = 256'h00008000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000001;
defparam prom_inst_3.INIT_RAM_32 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_33 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_34 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_35 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_36 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000800000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(prom_inst_2_dout[1]),
  .I1(prom_inst_3_dout[1]),
  .S0(dff_q_0)
);
endmodule //rom_4c
