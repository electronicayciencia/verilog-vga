//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Fri Dec 17 12:05:20 2021

module rom_font (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0010387CFEFEFE6C7EFFE7C3FFDBFF7E7E8199BD81A5817E0000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000183C3C18000038107CFEFE7C38103810D6FEFE387C380010387CFE7C3810;
defparam prom_inst_0.INIT_RAM_02 = 256'h78CCCCCC7D0F070FFFC399BDBD99C3FF003C664242663C00FFFFE7C3C3E7FFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'h18DB3CE7E73CDB18C0E66763637F637FE0F07030303F333F187E183C6666663C;
defparam prom_inst_0.INIT_RAM_04 = 256'h0066006666666666183C7E18187E3C1800020E3EFE3E0E020080E0F8FEF8E080;
defparam prom_inst_0.INIT_RAM_05 = 256'hFF183C7E187E3C18007E7E7E000000007C863C66663C613E001B1B1B7BDBDB7F;
defparam prom_inst_0.INIT_RAM_06 = 256'h00003060FE6030000000180CFE0C180000183C7E1818181800181818187E3C18;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000183C7EFFFF000000FFFF7E3C180000002466FF6624000000FEC0C0C00000;
defparam prom_inst_0.INIT_RAM_08 = 256'h006C6CFE6CFE6C6C000000000024666600180018183C3C180000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h00000000003018180076CCDC76386C3800C6663018CCC60000187C063C603E18;
defparam prom_inst_0.INIT_RAM_0A = 256'h000018187E1818000000663CFF3C66000030180C0C0C1830000C18303030180C;
defparam prom_inst_0.INIT_RAM_0B = 256'h0080C06030180C060018180000000000000000007E0000003018180000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h007CC6063C06C67C00FE66301C06C67C007E18181818381800386CC6D6C66C38;
defparam prom_inst_0.INIT_RAM_0D = 256'h00303030180CC6FE007CC6C6FCC06038007CC606FCC0C0FE001E0CFECC6C3C1C;
defparam prom_inst_0.INIT_RAM_0E = 256'h3018180000181800001818000018180000780C067EC6C67C007CC6C67CC6C67C;
defparam prom_inst_0.INIT_RAM_0F = 256'h00180018180CC67C006030180C18306000007E00007E000000060C1830180C06;
defparam prom_inst_0.INIT_RAM_10 = 256'h003C66C0C0C0663C00FC66667C6666FC00C6C6C6FEC66C380078C0DEDEDEC67C;
defparam prom_inst_0.INIT_RAM_11 = 256'h003A66CEC0C0663C00F06068786862FE00FE6268786862FE00F86C6666666CF8;
defparam prom_inst_0.INIT_RAM_12 = 256'h00E6666C786C66E60078CCCC0C0C0C1E003C18181818183C00C6C6C6FEC6C6C6;
defparam prom_inst_0.INIT_RAM_13 = 256'h007CC6C6C6C6C67C00C6C6CEDEF6E6C600C6C6D6FEFEEEC600FE6662606060F0;
defparam prom_inst_0.INIT_RAM_14 = 256'h003C660C1830663C00E6666C7C6666FC0E7CCEC6C6C6C67C00F060607C6666FC;
defparam prom_inst_0.INIT_RAM_15 = 256'h006CFED6D6C6C6C600386CC6C6C6C6C6007CC6C6C6C6C6C6003C1818185A7E7E;
defparam prom_inst_0.INIT_RAM_16 = 256'h003C30303030303C00FE6632188CC6FE003C18183C66666600C6C66C386CC6C6;
defparam prom_inst_0.INIT_RAM_17 = 256'hFF0000000000000000000000C66C3810003C0C0C0C0C0C3C0002060C183060C0;
defparam prom_inst_0.INIT_RAM_18 = 256'h007CC6C0C67C000000DC6666667C60E00076CC7C0C78000000000000000C1830;
defparam prom_inst_0.INIT_RAM_19 = 256'hF80C7CCCCC76000000F06060F860663C007CC0FEC67C00000076CCCCCC7C0C1C;
defparam prom_inst_0.INIT_RAM_1A = 256'h00E66C786C6660E03C66660606060006003C18181838001800E66666766C60E0;
defparam prom_inst_0.INIT_RAM_1B = 256'h007CC6C6C67C00000066666666DC000000D6D6D6FEEC0000003C181818181838;
defparam prom_inst_0.INIT_RAM_1C = 256'h00FC067CC07E000000F0606076DC00001E0C7CCCCC760000F0607C6666DC0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h006CFED6D6C6000000386CC6C6C600000076CCCCCCCC0000001C363030FC3030;
defparam prom_inst_0.INIT_RAM_1E = 256'h000E18187018180E007E32184C7E0000FC067EC6C6C6000000C66C386CC60000;
defparam prom_inst_0.INIT_RAM_1F = 256'h00FEC6C66C381000000000000000DC76007018180E1818700018181818181818;
defparam prom_inst_0.INIT_RAM_20 = 256'h0076CC7C0C78827C007CC0FEC67C180C0076CCCCCCCC00CC780C7CC6C0C0C67C;
defparam prom_inst_0.INIT_RAM_21 = 256'h380C7EC0C07E00000076CC7C0C7830300076CC7C0C7818300076CC7C0C7800C6;
defparam prom_inst_0.INIT_RAM_22 = 256'h003C181818380066007CC0FEC67C1830007CC0FEC67C00C6007CC0FEC67C827C;
defparam prom_inst_0.INIT_RAM_23 = 256'h00C6C6FEC67C6C3800C6C6FEC66C38C6003C181838001830003C18181838827C;
defparam prom_inst_0.INIT_RAM_24 = 256'h007CC6C6C67C827C00CECCCCFECC6C3E007ED87E187E000000FEC0F8C0FE3018;
defparam prom_inst_0.INIT_RAM_25 = 256'h0076CCCCCCCC30600076CCCCCC008478007CC6C6C67C1830007CC6C6C67C00C6;
defparam prom_inst_0.INIT_RAM_26 = 256'h18187EC0C07E1818007CC6C6C6C600C600386CC6C66C38C6FC067EC6C6C600C6;
defparam prom_inst_0.INIT_RAM_27 = 256'h0070D8183C181B0EC7C6CFC6FACCCCF818187E187E3C666600FC6660F0646C38;
defparam prom_inst_0.INIT_RAM_28 = 256'h0076CCCCCCCC3018007CC6C6C67C180C003C18183800180C0076CC7C0C783018;
defparam prom_inst_0.INIT_RAM_29 = 256'h00007C00386C6C3800007E003E6C6C3C00CEDEF6E600DC7600666666DC00DC76;
defparam prom_inst_0.INIT_RAM_2A = 256'h0FCC66337E6CE66300000606FE0000000000C0C0FE000000003E633018180018;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000CC663366CC0000003366CC66330000183C3C1818001806DF6A367A6CE663;
defparam prom_inst_0.INIT_RAM_2C = 256'h1818181818181818DD77DD77DD77DD77AA55AA55AA55AA558822882288228822;
defparam prom_inst_0.INIT_RAM_2D = 256'h363636FE00000000363636F636363636181818F818F81818181818F818181818;
defparam prom_inst_0.INIT_RAM_2E = 256'h363636F606FE00003636363636363636363636F606F63636181818F818F80000;
defparam prom_inst_0.INIT_RAM_2F = 256'h181818F800000000000000F818F81818000000FE36363636000000FE06F63636;
defparam prom_inst_0.INIT_RAM_30 = 256'h1818181F18181818181818FF00000000000000FF181818180000001F18181818;
defparam prom_inst_0.INIT_RAM_31 = 256'h36363637363636361818181F181F1818181818FF18181818000000FF00000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h363636F700FF0000000000FF00F7363636363637303F00000000003F30373636;
defparam prom_inst_0.INIT_RAM_33 = 256'h000000FF00FF1818363636F700F73636000000FF00FF00003636363730373636;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000003F36363636363636FF00000000181818FF00FF0000000000FF36363636;
defparam prom_inst_0.INIT_RAM_35 = 256'h363636FF363636363636363F000000001818181F181F00000000001F181F1818;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF1818181F00000000000000F818181818181818FF18FF1818;
defparam prom_inst_0.INIT_RAM_37 = 256'h00000000FFFFFFFF0F0F0F0F0F0F0F0FF0F0F0F0F0F0F0F0FFFFFFFF00000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h006C6C6C6CFE000000C0C0C0C0C0C6FE00CCC6CCD8CCCC780076DCC8DC760000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0018181818DC7600C07C6666666600000070D8D8D87E000000FEC6603060C6FE;
defparam prom_inst_0.INIT_RAM_3A = 256'h003C66663E0C180E00EE6C6CC6C66C3800386CC6FEC66C387E183C66663C187E;
defparam prom_inst_0.INIT_RAM_3B = 256'h00C6C6C6C6C67C00001E30607E60301EC0607EDBDB7E0C0600007EDBDB7E0000;
defparam prom_inst_0.INIT_RAM_3C = 256'h007E000C1830180C007E0030180C1830007E0018187E18180000FE00FE00FE00;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000DC7600DC7600000018007E00180070D8D8181818181818181818181B1B0E;
defparam prom_inst_0.INIT_RAM_3E = 256'h1C3C6CEC0C0C0C0F0000000018000000000000181800000000000000386C6C38;
defparam prom_inst_0.INIT_RAM_3F = 256'h000000000000000000003C3C3C3C00000000007C30180C78000000363636366C;

endmodule //rom_font
