//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Thu Dec 09 13:39:45 2021

module texture1_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h3B073B073B073AE7528A8410949294929492A514A514949294929492AD75AD75;
defparam prom_inst_0.INIT_RAM_01 = 256'hAD75AD758C7173AE632C632C841084108C71AD75AD75AD75AD75AD7584106B4D;
defparam prom_inst_0.INIT_RAM_02 = 256'h3B073B073B073AE73266738E738E8410841084307BEF84308430843094929492;
defparam prom_inst_0.INIT_RAM_03 = 256'h843084308C7173AE632C841084108C71AD75AD75AD75AD758C718C513B073B07;
defparam prom_inst_0.INIT_RAM_04 = 256'h4488448844883B073AE7528A738E738E738E8410843084108430843084309492;
defparam prom_inst_0.INIT_RAM_05 = 256'h8430843073AE73AE528A84108C71AD75AD75AD758C7184108C5184103B073B07;
defparam prom_inst_0.INIT_RAM_06 = 256'h3BA784304488448844883AE732664A49738E738E84107BEF843084107BEF7BEF;
defparam prom_inst_0.INIT_RAM_07 = 256'h73AE73AE3B673AC73266326684108C7184108C5184108C513BA73BA73B073BA7;
defparam prom_inst_0.INIT_RAM_08 = 256'h3BA7843094923BA744883BA73B0732663246738E738E7BEF738E738E7BEF8410;
defparam prom_inst_0.INIT_RAM_09 = 256'h73AE3AC73AC73B073B0732663266841084108C518C5184103BA742284A698410;
defparam prom_inst_0.INIT_RAM_0A = 256'h8430841094923BE73BE7AD75C6383B0732663246738E738E7BEF738E3AC73AC7;
defparam prom_inst_0.INIT_RAM_0B = 256'h3AC73AC73B077BEF7BEF3BA73266326684108410841084104228528A4A694A69;
defparam prom_inst_0.INIT_RAM_0C = 256'h8410841094923BA76B6D8430C6383B073B0732663246738E3B473AC73AC73B07;
defparam prom_inst_0.INIT_RAM_0D = 256'h3B073B077BEFB5963BE7A5343BA73266528A52AA528A326632663B0732664A69;
defparam prom_inst_0.INIT_RAM_0E = 256'h7BEF841084106B6D843084303BE7AD753B073B07326632463AC73AC76B4D3B07;
defparam prom_inst_0.INIT_RAM_0F = 256'h6B4D632CB596B596A5347BEF3BA73AE73266528A32663A873B073B073B073A87;
defparam prom_inst_0.INIT_RAM_10 = 256'h52AA8410841084107BEF84308430AD753B073AE7632C632CA534A534AD756B4D;
defparam prom_inst_0.INIT_RAM_11 = 256'h6B4D632CB596A5347BEFA5347BEF3AE73AE744289CD39CD39CD344483B073266;
defparam prom_inst_0.INIT_RAM_12 = 256'h3266328684108410841084108430AD753AE73AE773AEA534A534A534AD75A534;
defparam prom_inst_0.INIT_RAM_13 = 256'h3B073A87A5347BEF7BEF6B4D632C632C9CD344283B879CD34428A51444683B07;
defparam prom_inst_0.INIT_RAM_14 = 256'h3AC732667BEF841084308410843044883AE76B4D73AE73AE841073AEA534AD75;
defparam prom_inst_0.INIT_RAM_15 = 256'h3B073A873BA77BEF3246632C6B6D6B6D8C513BC744287BEFA514C61844684468;
defparam prom_inst_0.INIT_RAM_16 = 256'h3AC7326632668410841084303B873B873AE73B0773AE843084308410AD75A534;
defparam prom_inst_0.INIT_RAM_17 = 256'h6B4D3A87324632466B4D6B6D84108C5184103BA73B87A514C618C6183BE74468;
defparam prom_inst_0.INIT_RAM_18 = 256'h3AC73B073266528A84107BEF3B873AE73AE73B07841073AE843073AE8410A534;
defparam prom_inst_0.INIT_RAM_19 = 256'hAD756B4D3A8784108410841073AE73AE84103BA74448A5148C713BE73BE73286;
defparam prom_inst_0.INIT_RAM_1A = 256'h3AC73B073B073266528A528A32663AE73AE732663B67841073AE73AE8410A534;
defparam prom_inst_0.INIT_RAM_1B = 256'hBDF7AD753B273A87841073AE73AE84108410841044488C718C713B8732863AC7;
defparam prom_inst_0.INIT_RAM_1C = 256'h3B073AE73AE73B07AD75A534446844683AE73266322673AE841073AE73AE8430;
defparam prom_inst_0.INIT_RAM_1D = 256'hBDF7AD753B073A87841073AE841084108C518C518410528A328632863AC73AC7;
defparam prom_inst_0.INIT_RAM_1E = 256'h3B073AE73B073BA74488448844884468B5B63AE73266322673AE841084108430;
defparam prom_inst_0.INIT_RAM_1F = 256'h8430BDF7AD753B273A87841084108C518C5173AE32863AC73AC73AC73B073B07;
defparam prom_inst_0.INIT_RAM_20 = 256'hAD753AE73AE73B073B873BC74488AD75B5B6B5B63AE7326632263B67841073AE;
defparam prom_inst_0.INIT_RAM_21 = 256'h84308430BDF7448842283A87841052AA632C3AC73AC73BA73BA73BE73BE7AD75;
defparam prom_inst_0.INIT_RAM_22 = 256'hB5B644883AC7528A3B073BC73BC7B596AD75B5B6AD753AE73266322673AE8410;
defparam prom_inst_0.INIT_RAM_23 = 256'h73AE84308430BDF7448842283A873A873B073B073AC794923BE73BE7A534A534;
defparam prom_inst_0.INIT_RAM_24 = 256'hB5B63B47B5B6632C32663B473BC78C51B596B596AD75AD753AE732663AE773AE;
defparam prom_inst_0.INIT_RAM_25 = 256'h8430843084308430BDF7AD753A873B073B073AC7841084303BE73BE7A534B5B6;
defparam prom_inst_0.INIT_RAM_26 = 256'h738EAD75B5B6632C528A32663BC784108C518C51B596AD75A5143AE73AE773AE;
defparam prom_inst_0.INIT_RAM_27 = 256'h843073AE843084309CD3AD75632C3B073266843084303BE73BE73BE78C71B5B6;
defparam prom_inst_0.INIT_RAM_28 = 256'h8410B5B6AD75AD75632C4A693B8784107BEF8C517BEF7BEF4448A5143AE7528A;
defparam prom_inst_0.INIT_RAM_29 = 256'h73AE8430841084109CD33AE73AE73B073266528A843084303BA794928410B5B6;
defparam prom_inst_0.INIT_RAM_2A = 256'h841094929492AD75632C528A73AE841084107BEF7BEF444844486B4D6B4D528A;
defparam prom_inst_0.INIT_RAM_2B = 256'h73AE73AE73AE9CD33AE73AE73B073AE73B073266326684103BA7841084109492;
defparam prom_inst_0.INIT_RAM_2C = 256'h9492949294929492632C4A6973AE73AE7BEF7BEF442844283B073B073B073B07;
defparam prom_inst_0.INIT_RAM_2D = 256'h4228528A73AE3AE73AE73AE7446844683AE73AE7326632668410841094928410;
defparam prom_inst_0.INIT_RAM_2E = 256'h8410843094928430632C4A69528A73AE7BEF9CD33266528A6B4D7BEFB5B63B07;
defparam prom_inst_0.INIT_RAM_2F = 256'h52AA528A3AE73AE73AE7A53444684428AD753AE73AE7326632663BA794928410;
defparam prom_inst_0.INIT_RAM_30 = 256'h84108410841084103AC73AC7326632663266326632666B4D7BEF8C51B5B6B5B6;
defparam prom_inst_0.INIT_RAM_31 = 256'h52AA3AE73AE73AE784108C51442844289CF3AD75AD75AD7532663AA794928430;
defparam prom_inst_0.INIT_RAM_32 = 256'h841084106B6D3B273B073AC73AC732663266326632663BA78C51AD758C51B5B6;
defparam prom_inst_0.INIT_RAM_33 = 256'h3AA73AA73AE78C518410841084103BE79CF38C519CF3AD75AD7532663AA7632C;
defparam prom_inst_0.INIT_RAM_34 = 256'h326632663B073B07A534B59644684468B5963B07326632667BEF8C518C51B5B6;
defparam prom_inst_0.INIT_RAM_35 = 256'h326632668410841084108C519492841084109492A514A514C638C6383AA73266;
defparam prom_inst_0.INIT_RAM_36 = 256'h3B073B0784308430B5967BEF4468A534B596B5963B073AA77BEF7BEF8C51AD75;
defparam prom_inst_0.INIT_RAM_37 = 256'h528A528A84108C51841084108C518C51841084108C51A514A51444883B073B07;
defparam prom_inst_0.INIT_RAM_38 = 256'h3B077BEF84307BEF7BEF7BEF84308430A534A5343AA76B4D52AA7BEF7BEF8C51;
defparam prom_inst_0.INIT_RAM_39 = 256'h3AA73A87528A84108C5184108C5194928C5184108C51841084103B073B073B07;
defparam prom_inst_0.INIT_RAM_3A = 256'h3B073266843084307BEF84308430A534843032663AA752AA52AA52AA52AA52AA;
defparam prom_inst_0.INIT_RAM_3B = 256'h3AA73A873A87326684108C5194928C51841084108410632C3BA73B073B074488;
defparam prom_inst_0.INIT_RAM_3C = 256'h3B073266326632667BEF7BEF7BEF843032663AA7632CA514A514632C632C632C;
defparam prom_inst_0.INIT_RAM_3D = 256'h632C632C3AE73A8732663AA73AA73A873B073B07632C632C8410841044884488;
defparam prom_inst_0.INIT_RAM_3E = 256'h6B4D6B4D3B07326632463246324632463B07632CA514AD75AD75AD75A514A514;
defparam prom_inst_0.INIT_RAM_3F = 256'hAD758C71AD75632C3A873A873A873AA73B0784108C71AD75AD758C71AD754488;

endmodule //texture1_rom
