//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Thu Dec 16 21:23:22 2021

module charbuf_mono_64x64 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [11:0] ada;
input [7:0] din;
input [11:0] adb;

wire [27:0] sdpb_inst_0_dout_w;
wire [27:0] sdpb_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[27:0],dout[3:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 4;
defparam sdpb_inst_0.BIT_WIDTH_1 = 4;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h00000000000000000000000000000356F409849C3058404E10C79CC922031747;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h00000000000000000000000000000000A521705840E905C2D9704E1052970494;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h00000000000000000000000000000000000C356F7F2F2058405257093D9D0CC1;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h000000000000000000000000000000000000E5212745F03841205DFD058404E1;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000001EF309D0CB3F725221A058405217527;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h00000000000000000000000183413041840371C305840C5492041840371A0584;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h00000000000000000000000000000000E58304E10C4292025A25A05840521752;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000718341E3254E12035F9D5260584;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000A4E180E9042F730C102F603980BFF4058;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000D4875F305805F605DF8E1D058405D9407EFC;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h00000000000000000000000000000000C55240D54D54058409205804543520F3;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h000000000000000000000000000000000000E4875F840E905C987104FF4304E1;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h00000000000000000000000000000C4FF4305804875F8408396650E90310C4E1;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h00000000000000000000000000000C5D1C606F03595084970CB3F725221A0584;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000C4FF70957C5405840875F28407E9C6698705D13;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000015D13049031045C225204E1;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h000000000000000000000875F28404E10875F28404E101F740C5EF01F740C5EF;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h00000000000000000000000000001B31E3D25B39E304E570541C20C102F60584;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h000000000000000000000000000000415803490849704E10C41540490465C058;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000EB31207E980D5C1704E57058;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000FB3F725221A05840E91C305F840431804E17;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000019F20839D15209D0C3D2109D0F405DF3;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h00000000000000000000000000000007191CC13018FFCC1301914035FA21260F;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h00000000000000000000000000000000000000000E9FA03980E9045C42F83058;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h00000000000000000000000000000356F409849C3058404E10C79CC922031747;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h00000000000000000000000000000000A521705840E905C2D9704E1052970494;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h00000000000000000000000000000000000C356F7F2F2058405257093D9D0CC1;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h000000000000000000000000000000000000E5212745F03841205DFD058404E1;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[27:0],dout[7:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 4;
defparam sdpb_inst_1.BIT_WIDTH_1 = 4;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h2222222222222222222222222222276767276766726672666226666676276752;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h2222222222222222222222222222222236667266726626666662666267762664;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h2222222222222222222222222222222222227676667662667267672776662664;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h2222222222222222222222222222222222222666767762767672666626672664;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h2222222222222222222222222222222222667276226667766664266726767642;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h2222222222222222222222226676627667277666266722676627667277662665;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h2222222222222222222222222222222267672666226766267667426672676764;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h2222222222222222222222222222222222222226676677666642776667762665;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h2222222222222222222222222222222366662662676772667767276626667264;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h2222222222222222222222222222276676726626662666766626672666726664;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h2222222222222222222222222222222226677267767526672762662667767265;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h2222222222222222222222222222222222222766766726626666762666772664;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h2222222222222222222222222222226667726627667667267666726627622664;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h2222222222222222222222222222226666626627676267672266677666642665;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h2222222222222222222222222266672766677266726676767266666666726664;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h2222222222222222222222222222222222222222226666276276266667762664;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h2222222222222222222226676767266626676767266422677226642267722664;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h2222222222222222222222222222266667276666672766726666626677672665;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h2222222222222222222222222222226666277626767266622666627627666264;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h2222222222222222222222222222222222222222266662666676766627667264;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h2222222222222222222222222222366677666642667266667276672776626642;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h2222222222222222222222222222222227662676666627622767627626726664;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h2222222222222222222222222222222227666642266666642276627766667624;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h2222222222222222222222222222222222222222227662766266266677666264;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h2222222222222222222222222222276767276766726672666226666676276752;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h2222222222222222222222222222222236667266726626666662666267762664;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h2222222222222222222222222222222222227676667662667267672776662664;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h2222222222222222222222222222222222222666767762767672666626672664;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h2222222222222222222222222222222222222222222222222222222222222222;

endmodule //charbuf_mono_64x64
