//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Wed Dec 08 22:25:38 2021

module rom_led_off (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'hAD55A51494B28410630C10A20000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h000000000000000000000000000000000000000010A2630C841094B2A514AD55;
defparam prom_inst_0.INIT_RAM_04 = 256'hA534A534A534A534A5349CF37BCF294500000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000029457BCF9CF3A534A534A534A534A534;
defparam prom_inst_0.INIT_RAM_06 = 256'h9CF39CF3A514A514A514A514A5149CD3630C0000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000630C9CD3A514A514A514A514A5149CF39CF3;
defparam prom_inst_0.INIT_RAM_08 = 256'h834D8B8E8C1094B29CD39CF39CF39CF39CF37BCF086100000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000008617BCF9CF39CF39CF39CF39492843083AE834D834D;
defparam prom_inst_0.INIT_RAM_0A = 256'h78007800802081658B4D9C929CD39CD39CD39CD37BEF08610000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h000000000000000008617BEF9CD39CD39CD38C717BAE7A8A7904780078007800;
defparam prom_inst_0.INIT_RAM_0C = 256'h780080829186A249AACB9A8A93AE9CF394B294B294B273AE0000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h000000000000000073AE94B294B294B27BEF728A788278007800780078007800;
defparam prom_inst_0.INIT_RAM_0E = 256'h780080829145A228AAEBBBCFBBEF932C9CF394929492949252AA000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h00000000000052AA949294929492738E79E77800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_10 = 256'h78008041910499E7AACBBB8EC471C4B2934D9CF38C718C718C51210400000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000000021048C518C718C7173AE71C778007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_12 = 256'h7800802088E399A6AA8AB36DC430D514C4F393CF94B28C518C51632C00000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h00000000632C8C518C517BEF7228780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_14 = 256'h7800800088A29186A249B32CBBEFCCD3DDB6ABAEA4F38C518430841008610000;
defparam prom_inst_0.INIT_RAM_15 = 256'h000008618410843084306AEB7861780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_16 = 256'h7800780080619145A228AAEBBBCFCC92D575CD55938E9492841084104A490000;
defparam prom_inst_0.INIT_RAM_17 = 256'h00004A498410841073AE71E77800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_18 = 256'h780078008041910499E7AACBBB8EC471D534DDF781869CF37BEF7BEF630C0000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000630C7BEF7BEF632C78A27800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_1A = 256'h78007800780088A299A6A28AB34DC430D514DDB678009CB27BEF7BCF6B6D0000;
defparam prom_inst_0.INIT_RAM_1B = 256'h00006B6D7BCF7BCF628A78007800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_1C = 256'h780078007800780088E3A228B32CBBEFCCD3B41078009430841073AE738E0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000738E73AE73AE620878007800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_1E = 256'h78007800780078007800780089869A6992497800780093EF8410738E738E0000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000738E738E6B6D69E778007800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_20 = 256'h7800780078007800780078007800780078007800780093EF7BEF6B6D6B6D0000;
defparam prom_inst_0.INIT_RAM_21 = 256'h00006B6D6B6D6B4D61E778007800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_22 = 256'h7800780078007800780078007800780078007800780094107BCF6B4D6B4D0000;
defparam prom_inst_0.INIT_RAM_23 = 256'h00006B4D6B4D6B4D61E778007800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_24 = 256'h780078007800780078007800780078007800780078009C926B4D632C5AEB0000;
defparam prom_inst_0.INIT_RAM_25 = 256'h00005AEB632C632C5A4978007800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_26 = 256'h780078007800780078007800780078007800780081659492632C632C4A690000;
defparam prom_inst_0.INIT_RAM_27 = 256'h00004A69632C632C52AA78827800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_28 = 256'h78007800780078007800780078007800780078008B4D7BEF630C630C31A60000;
defparam prom_inst_0.INIT_RAM_29 = 256'h000031A6630C630C5ACB69A67800780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_2A = 256'h78007800780078007800780078007800780080E39471630C5AEB5ACB00200000;
defparam prom_inst_0.INIT_RAM_2B = 256'h000000205ACB5AEB5AEB52697841780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_2C = 256'h7800780078007800780078007800780078008B6D73AE5ACB5ACB39E700000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000000039E75ACB5ACB52AA69C7780078007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_2E = 256'h7800780078007800780078007800780082AA843052AA52AA528A108200000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h000000001082528A52AA52AA528A716578007800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_30 = 256'h7800780078007800780078007800828A841052AA528A528A2965000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000000002965528A528A528A528A71657800780078007800780078007800;
defparam prom_inst_0.INIT_RAM_32 = 256'h7800780078007800780078A2832C7BCF528A4A694A6939C70000000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h000000000000000039C74A694A694A69528A6A08786178007800780078007800;
defparam prom_inst_0.INIT_RAM_34 = 256'h78007800780079047AAA7BAE632C4A494A494A4939E700200000000000000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000000000000000002039E74A494A494A494A695A8A71E778C3780078007800;
defparam prom_inst_0.INIT_RAM_36 = 256'h72AA72CB734D6B6D5AEB4A4942284228422831A6000000000000000000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h00000000000000000000000031A642284228422842284A695ACB6ACB728A728A;
defparam prom_inst_0.INIT_RAM_38 = 256'h4A694A694208420842084208420839E721240000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000212439E7420842084208420842084A494A49;
defparam prom_inst_0.INIT_RAM_3A = 256'h39E739E739E739E739E739E72965084100000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h000000000000000000000000000000000841296539E739E739E739E739E739E7;
defparam prom_inst_0.INIT_RAM_3C = 256'h39C739C73186296518E300000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000018E32965318639C739C7;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //rom_led_off
