//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Thu Dec 09 13:43:50 2021

module texture0_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h94B294B294B294B29CF39492949294929CF39CF39CF3A5149CD39CD39CD39CF3;
defparam prom_inst_0.INIT_RAM_01 = 256'h630C630C8C718C718C718C718C718C719CD39CD39CD394B294B294B294B294B2;
defparam prom_inst_0.INIT_RAM_02 = 256'h8C718C718C719492949294928C5194929492949294B294B294B2949294B29CF3;
defparam prom_inst_0.INIT_RAM_03 = 256'h630C5AEB73AE8C518C518C518C519492949294928C718C718C718C718C718C71;
defparam prom_inst_0.INIT_RAM_04 = 256'h8C518C518C518C518C518C517BCF7BCF8C518C518C517BEF7BEF8C5194929CF3;
defparam prom_inst_0.INIT_RAM_05 = 256'h630C5AEB73AE73AE7BEF7BEF7BEF7BCF7BCF7BCF7BCF7BCF7BEF7BEF738E8C51;
defparam prom_inst_0.INIT_RAM_06 = 256'h8C517BEF7BEF7BEF8C517BCF7BCF7BCF7BCF7BCF8C518C518C518C5194929CF3;
defparam prom_inst_0.INIT_RAM_07 = 256'h5AEB5AEB6B4D73AE7BEF7BCF7BCF7BEF7BCF7BCF7BEF7BEF7BEF738E738E738E;
defparam prom_inst_0.INIT_RAM_08 = 256'h7BEF7BEF8C518C517BCF7BCF8C518C517BCF7BCF7BCF7BCF7BCF7BEF94929492;
defparam prom_inst_0.INIT_RAM_09 = 256'h5AEB5ACB6B4D738E738E738E7BEF7BEF7BEF7BEF7BEF7BEF8C518C518C517BEF;
defparam prom_inst_0.INIT_RAM_0A = 256'h7BCF7BEF7BEF7BCF7BCF7BEF8C518C518C518C517BCF7BCF7BCF7BCF8C519492;
defparam prom_inst_0.INIT_RAM_0B = 256'h5AEB5ACB6B4D738E738E738E738E7BEF7BEF7BEF8C518C518C517BEF7BEF7BCF;
defparam prom_inst_0.INIT_RAM_0C = 256'h7BCF7BCF7BCF7BCF7BEF7BEF7BEF7BEF7BEF8C517BEF7BEF738E738E8C5194B2;
defparam prom_inst_0.INIT_RAM_0D = 256'h5AEB5ACB6B6D738E8C518C51738E7BEF7BEF7BCF7BCF7BCF7BEF7BEF7BEF7BEF;
defparam prom_inst_0.INIT_RAM_0E = 256'h7BCF7BCF7BEF7BEF7BEF8C518C518C517BEF7BEF7BEF738E738E7BCF8C7194B2;
defparam prom_inst_0.INIT_RAM_0F = 256'h5AEB5ACB6B6D738E8C517BEF7BEF7BEF7BEF7BEF7BEF7BCF7BCF7BCF7BCF7BCF;
defparam prom_inst_0.INIT_RAM_10 = 256'h8C518C517BCF7BCF7BCF7BCF7BCF8C518C517BCF7BCF7BCF7BCF7BCF8C7194B2;
defparam prom_inst_0.INIT_RAM_11 = 256'h5AEB5ACB6B6D73AE8C518C517BEF738E738E738E8C517BEF7BEF7BEF7BEF8C51;
defparam prom_inst_0.INIT_RAM_12 = 256'h8C518C518C518C517BCF7BCF7BCF7BCF7BCF7BCF7BCF7BCF7BCF7BCF8C7194B2;
defparam prom_inst_0.INIT_RAM_13 = 256'h5AEB5ACB73AE73AE7BEF8C517BEF7BEF7BEF738E738E8C518C518C518C518C51;
defparam prom_inst_0.INIT_RAM_14 = 256'h8C517BEF738E738E738E738E7BEF7BEF7BCF7BCF7BEF7BEF7BEF7BCF8C7194B2;
defparam prom_inst_0.INIT_RAM_15 = 256'h5AEB5AEB73AE738E7BCF7BCF7BCF7BEF7BEF7BEF738E738E7BCF7BCF7BEF8C51;
defparam prom_inst_0.INIT_RAM_16 = 256'h7BEF7BEF7BEF7BEF738E738E738E7BEF7BEF7BEF7BCF7BCF7BCF7BCF8C718C71;
defparam prom_inst_0.INIT_RAM_17 = 256'h630C5AEB6B4D738E7BEF7BEF7BCF7BCF7BCF7BEF7BEF7BCF7BCF7BCF7BCF7BCF;
defparam prom_inst_0.INIT_RAM_18 = 256'h738E738E738E738E738E738E738E73AE73AE73AE7BCF73AE73AE73AE8C518C71;
defparam prom_inst_0.INIT_RAM_19 = 256'h630C5AEB6B4D738E73AE738E738E738E6B6D73AE73AE73AE73AE73AE73AE73AE;
defparam prom_inst_0.INIT_RAM_1A = 256'h6B6D6B6D6B6D6B6D6B6D6B6D73AE73AE73AE7BCF7BCF7BCF738E738E738E8C71;
defparam prom_inst_0.INIT_RAM_1B = 256'h5AEB5AEB6B4D73AE73AE73AE6B6D632C632C632C738E738E73AE73AE73AE6B6D;
defparam prom_inst_0.INIT_RAM_1C = 256'h52AA5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5AEB;
defparam prom_inst_0.INIT_RAM_1D = 256'h5AEB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5AEB5AEB5AEB5ACB5ACB5ACB52AA52AA;
defparam prom_inst_0.INIT_RAM_1E = 256'h5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB;
defparam prom_inst_0.INIT_RAM_1F = 256'h5AEB5AEB5AEB5AEB630C630C630C630C630C630C630C630C5AEB5AEB5AEB5ACB;
defparam prom_inst_0.INIT_RAM_20 = 256'h5AEB5AEB94B294B29CF39CF39CF39CF394B294B294B294B294B294B294B29CF3;
defparam prom_inst_0.INIT_RAM_21 = 256'h9CF39CF394929CF39CF39CD39CD38C718C718C719CD39CF39CF39CF3A534A534;
defparam prom_inst_0.INIT_RAM_22 = 256'h5AEB5ACB6B6D8C718C7194929492949294928C718C718C718C718C718C718C71;
defparam prom_inst_0.INIT_RAM_23 = 256'h94928C518C518C5194929492949294928C5194929492949294B29CD39CD3A534;
defparam prom_inst_0.INIT_RAM_24 = 256'h5AEB5ACB6B6D73AE7BEF7BEF738E738E7BCF7BCF7BEF7BEF7BEF7BEF7BCF7BCF;
defparam prom_inst_0.INIT_RAM_25 = 256'h7BCF7BCF7BEF7BEF7BCF7BCF7BCF7BCF7BEF7BEF8C518C518C518C518C71A534;
defparam prom_inst_0.INIT_RAM_26 = 256'h5AEB5ACB73AE73AE7BEF7BEF7BEF738E738E738E738E7BCF7BCF7BEF7BEF7BEF;
defparam prom_inst_0.INIT_RAM_27 = 256'h7BCF7BCF7BCF7BEF7BEF7BEF7BEF7BEF7BEF7BEF7BEF7BEF8C518C518C7194B2;
defparam prom_inst_0.INIT_RAM_28 = 256'h630C5ACB73AE7BCF8C518C517BCF7BCF7BCF738E7BCF7BCF8C518C517BCF7BEF;
defparam prom_inst_0.INIT_RAM_29 = 256'h7BEF7BCF7BCF7BCF8C518C518C517BEF7BEF8C518C517BEF7BEF7BEF8C7194B2;
defparam prom_inst_0.INIT_RAM_2A = 256'h630C5ACB73AE738E8C518C518C518C517BCF7BCF7BCF8C518C518C518C518C51;
defparam prom_inst_0.INIT_RAM_2B = 256'h7BEF7BEF8C518C518C518C517BEF7BEF7BEF7BEF7BEF8C518C518C518C7194B2;
defparam prom_inst_0.INIT_RAM_2C = 256'h5AEB5ACB6B6D738E7BEF7BEF7BEF7BEF8C518C518C517BEF7BEF8C517BEF7BEF;
defparam prom_inst_0.INIT_RAM_2D = 256'h8C518C518C517BEF7BEF7BEF7BEF7BEF738E738E738E7BEF8C517BEF8C719CF3;
defparam prom_inst_0.INIT_RAM_2E = 256'h5AEB5ACB6B6D738E7BEF7BEF8C518C518C517BEF7BEF7BEF7BEF7BEF7BEF7BCF;
defparam prom_inst_0.INIT_RAM_2F = 256'h7BCF7BCF7BEF7BEF7BEF7BCF7BCF7BCF7BEF738E738E738E738E8C5194929CF3;
defparam prom_inst_0.INIT_RAM_30 = 256'h5AEB5ACB6B6D6B6D7BCF7BCF7BEF8C518C518C517BCF7BCF7BCF7BCF7BCF7BCF;
defparam prom_inst_0.INIT_RAM_31 = 256'h7BCF7BCF7BCF7BCF7BCF7BCF7BEF7BEF7BEF7BEF7BEF7BCF7BCF7BCF8C719CF3;
defparam prom_inst_0.INIT_RAM_32 = 256'h5AEB5ACB6B4D6B6D7BEF7BEF7BCF7BCF8C517BEF7BEF7BEF7BCF7BCF7BEF7BEF;
defparam prom_inst_0.INIT_RAM_33 = 256'h7BEF7BCF7BCF7BCF7BCF7BCF7BCF7BCF7BEF8C518C517BEF7BEF7BCF8C7194B2;
defparam prom_inst_0.INIT_RAM_34 = 256'h630C5ACB6B4D6B6D738E738E7BCF7BCF7BCF7BCF7BEF7BEF7BEF7BEF738E738E;
defparam prom_inst_0.INIT_RAM_35 = 256'h738E738E8C518C518C517BCF7BCF8C518C517BEF7BEF7BEF8C518C518C7194B2;
defparam prom_inst_0.INIT_RAM_36 = 256'h630C5AEB6B4D6B6D738E738E738E738E7BCF7BEF7BCF7BCF7BEF7BEF7BEF7BEF;
defparam prom_inst_0.INIT_RAM_37 = 256'h738E738E738E8C517BCF7BCF8C518C517BEF7BEF8C518C518C518C518C719492;
defparam prom_inst_0.INIT_RAM_38 = 256'h630C5AEB6B4D6B6D7BCF738E738E738E738E738E738E738E6B6D6B6D6B6D6B6D;
defparam prom_inst_0.INIT_RAM_39 = 256'h6B6D6B6D6B6D738E738E738E738E738E73AE7BCF7BCF7BCF738E738E8C718C51;
defparam prom_inst_0.INIT_RAM_3A = 256'h630C5ACB6B4D7BCF7BCF7BCF6B6D6B4D6B4D6B4D6B6D6B6D6B6D6B4D6B4D6B4D;
defparam prom_inst_0.INIT_RAM_3B = 256'h6B4D6B4D6B4D6B4D6B6D6B6D6B6D738E738E738E73AE73AE73AE6B6D6B6D8C51;
defparam prom_inst_0.INIT_RAM_3C = 256'h5AEB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB;
defparam prom_inst_0.INIT_RAM_3D = 256'h5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5ACB5AEB5ACB5ACB5ACB5ACB5AEB;
defparam prom_inst_0.INIT_RAM_3E = 256'h5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB630C630C630C5AEB;
defparam prom_inst_0.INIT_RAM_3F = 256'h5AEB5AEB5AEB5AEB5AEB5AEB5AEB5AEB630C630C630C630C5AEB5AEB5AEB5AEB;

endmodule //texture0_rom
