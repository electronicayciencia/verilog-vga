//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.03
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Thu Nov 02 22:09:34 2023

module charbuf_color_64x32 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [10:0] ada;
input [15:0] din;
input [10:0] adb;

wire [23:0] sdpb_inst_0_dout_w;
wire [23:0] sdpb_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[23:0],dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 8;
defparam sdpb_inst_0.BIT_WIDTH_1 = 8;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h093927D5A43F2C1B6685C232D51E21C6E422A56802490E4BE5183374F2C1B2AE;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h0000000013A2B2A3F97A63DE28276675AA67B4661AF96953E5E5E5687A6DD605;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hB9D60E7D6B457EE9B6BA23B3AB0B00EA30B72487E1EC1E9310E800C01B8D3655;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h00000000092EDC32FFBBDB99775844AC193CB05261138B68B91C9B53093FE1E8;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h5E10AFCA717C148B584652B2B8A5B78927FA2162B6AA2F2B253D4D3775C373A7;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h00000000D40EF8954422A1F620D02CC16360C3BE66A7028D00F78881E803BB36;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hF01FD2A8A374C9CFDAE90C309E1A1B7517559FB5572BEBFC538D0030F937AC64;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h00000000C3A2FB455AEEF4ABB394C1B2FFA8AD293871956ABB33732B6F231C62;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h14FC3F963C0AE97F567BED3B1F29C5A7199613F290538B28241F64C7FA7C288F;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h000000002DF4941C4FB96229344BF9962FB04928C6C34CBBF6FA09C7444C4368;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h3D9CBF0AEF7FAF65BF0CBF56C8811170EC37C8023700626CBE03B302B94A1BC0;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h000000004B3A68CF0FA8C7165D83A42744A08B6B13350CEEAC2BBC75B340B1D3;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h0FABF31221D7EA0EA38595ACAAA443EF3A7B4185C9D7D25F77AF28D592C25408;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h00000000E5281A5B9E4536D6EF455D55B62943F9791A60517E8BAE60F3AD2994;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h527111CF57ABAEB354C75B254DB0ECE74A8651EF95B80B934883180215566F37;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h000000001DC4D6CD97CD243AA59F8298F9A3CEA0C3DC7F4E3082753A1A7DDE11;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hE096DBD685A4F8A64EE42FD7B76E5EE9E5F2A08504D9986DAEFDA42763F2D965;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h00000000C2AEFEBA23DE106419C6EF577275F5BF5E5ABA3F2957EA7D8EE7928B;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h54939D9994F94CC281C3C77595433F291C28CCAF650762C80DCF2B94AE1D08D0;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h00000000E343E39E25F55047A185E7BAE1C54E81136D58520D3D87D642268A06;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hBD930FBEE50535F9AC5E3B7A90394AAF1C75C27E646D88C322D5F2484D3C35EE;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h000000007E60E439333F5B362B902DEA91073D43AB5DB7631B4274F376BC6856;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h4B9EC83F166ECCE2C929B8A047B71E45DA9F0305860D8D7CDC9956ADEAF54B81;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h0000000079C6A4E873632C17A0DCE7CE0A487930BD1CFC4995CD39254C94E091;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hE40A64EC708F6EBFC606590117A10AA6099A0165BD49A0D13F85C36B895F4A3F;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h00000000A8635B1BC0C5644A03CAE50227BC38F0B09D3CAC39AE06AF1732A8C4;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h76CA5D5DAE85561A1A42027F363BCF09C64A6CA782F1AE44033FD54F729B70DB;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h00000000E4EABE543CAC8CC1B7EAEA60DBBFD1510115C9F689EA5C9541AD94A5;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h4A7BA5F6E426F78A019176BAF1A2D1510F1C7720D9DF1D95D3AC3F4D98B8C70B;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h000000008B99BABCB43184E32D3A6A787890F469393F9A3CD745686258F85F8E;
defparam sdpb_inst_0.INIT_RAM_1E = 256'hA1682B4290AD519EF0982227B899D348AE0BD61F91FF7157C2607F0500C0795C;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h00000000082B775A1EAA908269F9490418C4997CE37BCB69338B027DDCE7EF0B;
defparam sdpb_inst_0.INIT_RAM_20 = 256'hDB265635B85990060E25463B2875A94BCB091DDDFF5710E2C7A676ED6F8AC926;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h0000000081B2ECBC3F757850CC5A3430011471E36B252938594BD504584CF1CC;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[23:0],dout[15:8]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:8]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 8;
defparam sdpb_inst_1.BIT_WIDTH_1 = 8;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h56DF72D0FF81461082EA6AD0BE600E676296AF6E1C822DE7DB7C45CE36A42303;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h000000001BAD519CBA0913D1556F49B0642F8C1D053BB1648AF759C783FEBF31;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h3F0D02143871AEFD37E787C2F63EE8D922FFE8148E54D6473CEDA7913563327C;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h00000000AB5A74B8ADCA08780B0D08A266592D2B28B4623097DE4BB0E3EC3930;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h46EC8613DA9F41B96A52507284D0D6F7E8ACA9015A6CC444AE4CBFE2B010D2CC;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h00000000B86C2F6D86A928897A1F9AB504DB895639BB135A200B077DD61ADE7D;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h2825B0BA63C030DEDBC4C5F72DD86FE67828CA7F58579D8B5C8AE9AA0A794603;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h00000000CEC14DF1C6B704F28EDE6A9271298F00677BF8D4B18C58FA2C031AD4;
defparam sdpb_inst_1.INIT_RAM_08 = 256'hDA6489E88547641D2D14B7CC87E607F39371F24DE00825E5B8871736DB455DC9;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h000000008F981A278CD0B5946BB354185339B463A9AF223A458EB26215A3DAAD;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h00440656278D58093CF324221F15D8358FCA8F58F954C647BAD46775F04BF542;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h00000000A6FC3814CFEF427122F3F07E51B45AA77BBBE136E797F8343B266FBA;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h9599AC1E03DD45787A68DE4747F71478F36C14363B4EC2B3BC0D09D0C2264B3E;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h000000004A57A010862C0893D91122A9DCCFC9608F6CCC1CD19FF1FAA4D5673D;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h874C990E253DE64E8F37BB869E31F47E0CCD1808FD4AC32B8BFC5160D4881704;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h00000000C89FD2DBC518E76D0DAACBBFFAD5F819C5BF366C371620DA473DE668;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hA8528B009893C2D8E736C07174CADC7C345CEC3802E65D08E971274498B0F4C7;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h00000000123F10CE5E1824108724CDD939789C4F2E4ADCB1E322C33CC803A13F;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hBB38B5D807684C3DB5411394AF53CAD282A6FB6EDF1BDF6A92A9AE00D8128DE6;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h000000006596E7B1A080EDE622A346C87C07C3B75B877BBD8296688A76D143AD;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h8F6A3C36E87C9A6FB693559776AB5C201CD1B6AA97EE0380B7EB911AF55B45AD;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h000000005D642487A9598CC86B27F8BFD84612ED4C55BB31807E7E0B227FF339;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h4105DBF0864DA6C098D9619F5BA63523E80AD5973D31FB22E5992C5EDA1D4CB8;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h0000000033258E37F3A9100EF6F14F4A28C022327B534E54141626A6AC66F57A;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h7BD3BB221FB5DF04AB197BC6AA9E342403B2EE162BE3A15B05B67F7E19C6CE45;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h000000000105814A6BB71460475544F61FD091AA949465CF743C92A4DAC9F504;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h367A56F718BF332C8672A1620F253F7E84B1CE959CDD56FAC3F7B86393093F86;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h0000000058615D06CF3B9C7C6D9B72D54CAE88247E8699C1A11CDD8E405B1A05;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hC5F738B12E7A8F801372002128DBE6854794E7B1B47DEE9DA6FE18714D713E5A;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h00000000CDAE511A261FE00778F18C1446F1D43804C40F66B952F088C6161634;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h49495AE925B9A9AA60FB2AE2AB1D3BEE7E374716A5A236A39252CA2825CE7049;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h00000000D08B5882007E0C1D699D1816677D37CE6B503568C7590E3C63073252;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h51FDEB912F11AF5B90062D60BB0BC53E8F868C9501E54FFF96F68340A0A53194;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h0000000057842E7636BC5E7D1217117EDE8B7C223BBCBA7D80A3B40044B75421;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //charbuf_color_64x32
